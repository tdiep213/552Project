/*
   CS/ECE 552 Spring '22
  
   Filename        : execute.v
   Description     : This is the overall module for the execute stage of the processor.
*/
`default_nettype none
module execute (/* TODO: Add appropriate inputs/outputs for your execute stage here*/);

   // TODO: Your code here
   
endmodule
`default_nettype wire
