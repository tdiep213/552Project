//Arithmetic module
module alu();
endmodule