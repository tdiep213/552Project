    /*
    CS/ECE 552 Spring '22

    Filename        : fetch.v
    Description     : This is the module for the branch and jump component of the processor
    */
`default_nettype none
    //Branch + Jump calculation
module brancher (BJAddr, RetAddr, PC, Imm, RegVal);

// Move over anything extra from PC

endmodule
`default_nettype wire