/*
   CS/ECE 552 Spring '22
  
   Filename        : fetch.v
   Description     : This is the module for the overall fetch stage of the processor.
*/
`default_nettype none
module fetch (/* TODO: Add appropriate inputs/outputs for your fetch stage here*/);

   // TODO: Your code here
   
endmodule
`default_nettype wire
