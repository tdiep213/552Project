module dm_fsm();
endmodule